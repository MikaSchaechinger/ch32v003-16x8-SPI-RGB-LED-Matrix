module Address_Generator #(
    parameter int ADDRESS_BITS = 8
) (
    input  logic                          I_rst_n,
    input  logic                          I_address_up,
    input  logic                          I_address_reset,
    
    output logic [ADDRESS_BITS-1:0]       O_address
);




endmodule